//the files is the demod module files
