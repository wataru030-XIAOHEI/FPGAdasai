module filter (
    
);

endmodule //filter