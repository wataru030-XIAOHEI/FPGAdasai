//the files is the ammod module file
